library verilog;
use verilog.vl_types.all;
entity t_transmitter is
end t_transmitter;

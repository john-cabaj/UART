library verilog;
use verilog.vl_types.all;
entity t_bus_interface is
end t_bus_interface;

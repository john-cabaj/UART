library verilog;
use verilog.vl_types.all;
entity t_baud_generator is
end t_baud_generator;

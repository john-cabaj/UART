library verilog;
use verilog.vl_types.all;
entity t_top_level_full is
end t_top_level_full;

library verilog;
use verilog.vl_types.all;
entity t_receiver is
end t_receiver;
